library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity comparateur is 
  port(
    A,B:in std_logic;
    S1,S2,S3: out std_logic);
end comparateur;

architecture behavioral of comparateur is
begin 
S1<='1' when (A<B) else '0';
S2<='1' when (A=B) else '0';
S3<='1' when (A>B) else '0';
end behavioral;
             