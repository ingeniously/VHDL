library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity Counting_Transcoder is 
  port(
    H: in std_logic;
    O: out std_logic_vector(6 downto 0));
end Counting_Transcoder;

architecture behavioral of Counting_Transcoder is
 
signal C: std_logic_vector(3 downto 0);

  
   component Horloge 
     port(
         H:in std_logic;
         S: out std_logic_vector(4 downto 1):="0000");
   end component;

  component Transcoder 
  port(
    E: in std_logic_vector(3 downto 0);
    S: out std_logic_vector(6 downto 0));
  end component;

begin
u1: Horloge port map (H,C);
u2: Transcoder port map (C,O);
end behavioral;